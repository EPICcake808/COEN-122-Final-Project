module assembly_code();
  assign instr[0] = 32'b01110001000001000001000000000000 //SUB x4, x4, x4
  assign instr[1] = 32'b01000001010000100000110000000000 //ADD x5, x2, x3
  assign instr[2] = 32'b11110010010000000000010000000001 //SVPC x9, 1
  assign instr[3] = 32'b11100001100000100000000000000000 //LD x6, x2
  assign instr[4] = 32'b00000000000000000000000000000000 //NOP
  assign instr[5] = 32'b00000000000000000000000000000000 //NOP
  assign instr[6] = 32'b01000001000001000001100000000000 //ADD x4, x4, x6
  assign instr[7] = 32'b01010000100000100000010000000000 //INC x2, x2, 1
  assign instr[8] = 32'b00000000000000000000000000000000 //NOP
  assign instr[9] = 32'b00000000000000000000000000000000 //NOP
  assign instr[10] = 32'b01110010000000100001010000000000 //SUB x8, x2, x5
  assign instr[11] = 32'b10110000000010010000000000000000 //BRN x9
  
endmodule
